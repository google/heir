// RUN: run_verilog \
// RUN:  --verilog_module %s \
// RUN:  --input='arg1=0' \
// RUN:  --input='arg1=128' \
// RUN:  --input='arg1=-64' \
// RUN:  --input='arg1=64' \
// RUN:  > %t
// RUN: FileCheck %s < %t

// CHECK: b'\x04'
// CHECK-NEXT: b'\x04'
// CHECK-NEXT: b'\x7e'
// CHECK-NEXT: b'\x82'
module main(
  input wire signed [7:0] arg1,
  output wire signed [7:0] _out_
);
  wire signed [31:0] v2;
  wire signed [31:0] v3;
  wire signed [63:0] v4;
  wire signed [63:0] v5;
  wire signed [31:0] v6;
  wire signed [7:0] v7;
  wire signed [7:0] v8;
  wire signed [31:0] v9;
  wire signed [63:0] v10;
  wire signed [63:0] v11;
  wire signed [63:0] v12;
  wire signed [63:0] v13;
  wire signed [63:0] v14;
  wire signed [63:0] v15;
  wire signed [63:0] v16;
  wire signed [63:0] v17;
  wire signed [63:0] v18;
  wire signed [31:0] v19;
  wire signed [31:0] v20;
  wire signed [31:0] v21;
  wire signed [31:0] v22;
  wire signed [31:0] v23;
  wire signed [31:0] v24;
  wire signed [31:0] v25;
  wire signed [31:0] v26;
  wire signed [31:0] v27;
  wire signed [31:0] v28;
  wire signed [31:0] v29;
  wire signed [31:0] v30;
  wire signed [31:0] v31;
  wire signed [31:0] v32;
  wire signed [31:0] v33;
  wire signed [31:0] v34;
  wire signed [31:0] v35;
  wire signed [31:0] v36;
  wire signed [31:0] v37;
  wire signed [31:0] v38;
  wire signed [31:0] v39;
  wire signed [31:0] v40;
  wire signed [31:0] v41;
  wire signed [31:0] v42;
  wire signed [31:0] v43;
  wire signed [31:0] v44;
  wire signed [31:0] v45;
  wire signed [31:0] v46;
  wire signed [31:0] v47;
  wire signed [31:0] v48;
  wire signed [31:0] v49;
  wire signed [31:0] v50;
  wire signed [31:0] v51;
  wire signed [31:0] v52;
  wire signed [31:0] v53;
  wire signed [31:0] v54;
  wire signed [31:0] v55;
  wire signed [31:0] v56;
  wire signed [31:0] v57;
  wire signed [31:0] v58;
  wire signed [31:0] v59;
  wire signed [31:0] v60;
  wire signed [31:0] v61;
  wire signed [31:0] v62;
  wire signed [31:0] v63;
  wire signed [31:0] v64;
  wire signed [31:0] v65;
  wire signed [31:0] v66;
  wire signed [31:0] v67;
  wire signed [31:0] v68;
  wire signed [31:0] v69;
  wire signed [31:0] v70;
  wire signed [31:0] v71;
  wire signed [31:0] v72;
  wire signed [31:0] v73;
  wire signed [31:0] v74;
  wire signed [31:0] v75;
  wire signed [31:0] v76;
  wire signed [31:0] v77;
  wire signed [31:0] v78;
  wire signed [31:0] v79;
  wire signed [31:0] v80;
  wire signed [31:0] v81;
  wire signed [31:0] v82;
  wire signed [31:0] v83;
  wire signed [31:0] v84;
  wire signed [31:0] v85;
  wire signed [31:0] v86;
  wire signed [31:0] v87;
  wire signed [31:0] v88;
  wire signed [31:0] v89;
  wire signed [31:0] v90;
  wire signed [31:0] v91;
  wire signed [31:0] v92;
  wire signed [31:0] v93;
  wire signed [31:0] v94;
  wire signed [31:0] v95;
  wire signed [31:0] v96;
  wire signed [31:0] v97;
  wire signed [31:0] v98;
  wire signed [31:0] v99;
  wire signed [31:0] v100;
  wire signed [31:0] v101;
  wire signed [31:0] v102;
  wire signed [31:0] v103;
  wire signed [31:0] v104;
  wire signed [31:0] v105;
  wire signed [31:0] v106;
  wire signed [31:0] v107;
  wire signed [31:0] v108;
  wire signed [31:0] v109;
  wire signed [31:0] v110;
  wire signed [31:0] v111;
  wire signed [31:0] v112;
  wire signed [31:0] v113;
  wire signed [31:0] v114;
  wire signed [31:0] v115;
  wire signed [31:0] v116;
  wire signed [31:0] v117;
  wire signed [31:0] v118;
  wire signed [31:0] v119;
  wire signed [31:0] v120;
  wire signed [31:0] v121;
  wire signed [31:0] v122;
  wire signed [31:0] v123;
  wire signed [31:0] v124;
  wire signed [31:0] v125;
  wire signed [31:0] v126;
  wire signed [31:0] v127;
  wire signed [31:0] v128;
  wire signed [31:0] v129;
  wire signed [31:0] v130;
  wire signed [31:0] v131;
  wire signed [31:0] v132;
  wire signed [31:0] v133;
  wire signed [31:0] v134;
  wire signed [31:0] v135;
  wire signed [31:0] v136;
  wire signed [31:0] v137;
  wire signed [31:0] v138;
  wire signed [31:0] v139;
  wire signed [31:0] v140;
  wire signed [31:0] v141;
  wire signed [31:0] v142;
  wire signed [31:0] v143;
  wire signed [31:0] v144;
  wire signed [31:0] v145;
  wire signed [31:0] v146;
  wire signed [31:0] v147;
  wire signed [31:0] v148;
  wire signed [31:0] v149;
  wire signed [31:0] v150;
  wire signed [31:0] v151;
  wire signed [31:0] v152;
  wire signed [31:0] v153;
  wire signed [31:0] v154;
  wire signed [31:0] v155;
  wire signed [31:0] v156;
  wire signed [31:0] v157;
  wire signed [31:0] v158;
  wire signed [31:0] v159;
  wire signed [31:0] v160;
  wire signed [31:0] v161;
  wire signed [31:0] v162;
  wire signed [31:0] v163;
  wire signed [31:0] v164;
  wire signed [31:0] v165;
  wire signed [31:0] v166;
  wire signed [31:0] v167;
  wire signed [31:0] v168;
  wire signed [31:0] v169;
  wire signed [31:0] v170;
  wire signed [31:0] v171;
  wire signed [31:0] v172;
  wire signed [31:0] v173;
  wire signed [63:0] v174;
  wire signed [63:0] v175;
  wire signed [63:0] v176;
  wire v177;
  wire signed [63:0] v178;
  wire signed [63:0] v179;
  wire signed [63:0] v180;
  wire signed [31:0] v181;
  wire signed [31:0] v182;
  wire v183;
  wire signed [31:0] v184;
  wire v185;
  wire signed [31:0] v186;
  wire signed [7:0] v187;
  wire signed [63:0] v188;
  wire signed [63:0] v189;
  wire signed [63:0] v190;
  wire v191;
  wire signed [63:0] v192;
  wire signed [63:0] v193;
  wire signed [63:0] v194;
  wire signed [31:0] v195;
  wire signed [31:0] v196;
  wire v197;
  wire signed [31:0] v198;
  wire v199;
  wire signed [31:0] v200;
  wire signed [7:0] v201;
  wire signed [63:0] v202;
  wire signed [63:0] v203;
  wire signed [63:0] v204;
  wire v205;
  wire signed [63:0] v206;
  wire signed [63:0] v207;
  wire signed [63:0] v208;
  wire signed [31:0] v209;
  wire signed [31:0] v210;
  wire v211;
  wire signed [31:0] v212;
  wire v213;
  wire signed [31:0] v214;
  wire signed [7:0] v215;
  wire signed [63:0] v216;
  wire signed [63:0] v217;
  wire signed [63:0] v218;
  wire v219;
  wire signed [63:0] v220;
  wire signed [63:0] v221;
  wire signed [63:0] v222;
  wire signed [31:0] v223;
  wire signed [31:0] v224;
  wire v225;
  wire signed [31:0] v226;
  wire v227;
  wire signed [31:0] v228;
  wire signed [7:0] v229;
  wire signed [63:0] v230;
  wire signed [63:0] v231;
  wire signed [63:0] v232;
  wire v233;
  wire signed [63:0] v234;
  wire signed [63:0] v235;
  wire signed [63:0] v236;
  wire signed [31:0] v237;
  wire signed [31:0] v238;
  wire v239;
  wire signed [31:0] v240;
  wire v241;
  wire signed [31:0] v242;
  wire signed [7:0] v243;
  wire signed [63:0] v244;
  wire signed [63:0] v245;
  wire signed [63:0] v246;
  wire v247;
  wire signed [63:0] v248;
  wire signed [63:0] v249;
  wire signed [63:0] v250;
  wire signed [31:0] v251;
  wire signed [31:0] v252;
  wire v253;
  wire signed [31:0] v254;
  wire v255;
  wire signed [31:0] v256;
  wire signed [7:0] v257;
  wire signed [63:0] v258;
  wire signed [63:0] v259;
  wire signed [63:0] v260;
  wire v261;
  wire signed [63:0] v262;
  wire signed [63:0] v263;
  wire signed [63:0] v264;
  wire signed [31:0] v265;
  wire signed [31:0] v266;
  wire v267;
  wire signed [31:0] v268;
  wire v269;
  wire signed [31:0] v270;
  wire signed [7:0] v271;
  wire signed [63:0] v272;
  wire signed [63:0] v273;
  wire signed [63:0] v274;
  wire v275;
  wire signed [63:0] v276;
  wire signed [63:0] v277;
  wire signed [63:0] v278;
  wire signed [31:0] v279;
  wire signed [31:0] v280;
  wire v281;
  wire signed [31:0] v282;
  wire v283;
  wire signed [31:0] v284;
  wire signed [7:0] v285;
  wire signed [63:0] v286;
  wire signed [63:0] v287;
  wire signed [63:0] v288;
  wire v289;
  wire signed [63:0] v290;
  wire signed [63:0] v291;
  wire signed [63:0] v292;
  wire signed [31:0] v293;
  wire signed [31:0] v294;
  wire v295;
  wire signed [31:0] v296;
  wire v297;
  wire signed [31:0] v298;
  wire signed [7:0] v299;
  wire signed [63:0] v300;
  wire signed [63:0] v301;
  wire signed [63:0] v302;
  wire v303;
  wire signed [63:0] v304;
  wire signed [63:0] v305;
  wire signed [63:0] v306;
  wire signed [31:0] v307;
  wire signed [31:0] v308;
  wire v309;
  wire signed [31:0] v310;
  wire v311;
  wire signed [31:0] v312;
  wire signed [7:0] v313;
  wire signed [63:0] v314;
  wire signed [63:0] v315;
  wire signed [63:0] v316;
  wire v317;
  wire signed [63:0] v318;
  wire signed [63:0] v319;
  wire signed [63:0] v320;
  wire signed [31:0] v321;
  wire signed [31:0] v322;
  wire v323;
  wire signed [31:0] v324;
  wire v325;
  wire signed [31:0] v326;
  wire signed [7:0] v327;
  wire signed [63:0] v328;
  wire signed [63:0] v329;
  wire signed [63:0] v330;
  wire v331;
  wire signed [63:0] v332;
  wire signed [63:0] v333;
  wire signed [63:0] v334;
  wire signed [31:0] v335;
  wire signed [31:0] v336;
  wire v337;
  wire signed [31:0] v338;
  wire v339;
  wire signed [31:0] v340;
  wire signed [7:0] v341;
  wire signed [63:0] v342;
  wire signed [63:0] v343;
  wire signed [63:0] v344;
  wire v345;
  wire signed [63:0] v346;
  wire signed [63:0] v347;
  wire signed [63:0] v348;
  wire signed [31:0] v349;
  wire signed [31:0] v350;
  wire v351;
  wire signed [31:0] v352;
  wire v353;
  wire signed [31:0] v354;
  wire signed [7:0] v355;
  wire signed [63:0] v356;
  wire signed [63:0] v357;
  wire signed [63:0] v358;
  wire v359;
  wire signed [63:0] v360;
  wire signed [63:0] v361;
  wire signed [63:0] v362;
  wire signed [31:0] v363;
  wire signed [31:0] v364;
  wire v365;
  wire signed [31:0] v366;
  wire v367;
  wire signed [31:0] v368;
  wire signed [7:0] v369;
  wire signed [63:0] v370;
  wire signed [63:0] v371;
  wire signed [63:0] v372;
  wire v373;
  wire signed [63:0] v374;
  wire signed [63:0] v375;
  wire signed [63:0] v376;
  wire signed [31:0] v377;
  wire signed [31:0] v378;
  wire v379;
  wire signed [31:0] v380;
  wire v381;
  wire signed [31:0] v382;
  wire signed [7:0] v383;
  wire signed [63:0] v384;
  wire signed [63:0] v385;
  wire signed [63:0] v386;
  wire v387;
  wire signed [63:0] v388;
  wire signed [63:0] v389;
  wire signed [63:0] v390;
  wire signed [31:0] v391;
  wire signed [31:0] v392;
  wire v393;
  wire signed [31:0] v394;
  wire v395;
  wire signed [31:0] v396;
  wire signed [7:0] v397;
  wire v398;
  wire signed [7:0] v399;
  wire v400;
  wire signed [7:0] v401;
  wire v402;
  wire signed [7:0] v403;
  wire v404;
  wire signed [7:0] v405;
  wire v406;
  wire signed [7:0] v407;
  wire v408;
  wire signed [7:0] v409;
  wire v410;
  wire signed [7:0] v411;
  wire v412;
  wire signed [7:0] v413;
  wire v414;
  wire signed [7:0] v415;
  wire v416;
  wire signed [7:0] v417;
  wire v418;
  wire signed [7:0] v419;
  wire v420;
  wire signed [7:0] v421;
  wire v422;
  wire signed [7:0] v423;
  wire v424;
  wire signed [7:0] v425;
  wire v426;
  wire signed [7:0] v427;
  wire v428;
  wire signed [7:0] v429;
  wire v430;
  wire signed [7:0] v431;
  wire v432;
  wire signed [7:0] v433;
  wire v434;
  wire signed [7:0] v435;
  wire v436;
  wire signed [7:0] v437;
  wire v438;
  wire signed [7:0] v439;
  wire v440;
  wire signed [7:0] v441;
  wire v442;
  wire signed [7:0] v443;
  wire v444;
  wire signed [7:0] v445;
  wire v446;
  wire signed [7:0] v447;
  wire v448;
  wire signed [7:0] v449;
  wire v450;
  wire signed [7:0] v451;
  wire v452;
  wire signed [7:0] v453;
  wire v454;
  wire signed [7:0] v455;
  wire v456;
  wire signed [7:0] v457;
  wire v458;
  wire signed [7:0] v459;
  wire v460;
  wire signed [7:0] v461;
  wire signed [31:0] v462;
  wire signed [31:0] v463;
  wire signed [31:0] v464;
  wire signed [31:0] v465;
  wire signed [31:0] v466;
  wire signed [31:0] v467;
  wire signed [31:0] v468;
  wire signed [31:0] v469;
  wire signed [31:0] v470;
  wire signed [31:0] v471;
  wire signed [31:0] v472;
  wire signed [31:0] v473;
  wire signed [31:0] v474;
  wire signed [31:0] v475;
  wire signed [31:0] v476;
  wire signed [31:0] v477;
  wire signed [31:0] v478;
  wire signed [31:0] v479;
  wire signed [31:0] v480;
  wire signed [31:0] v481;
  wire signed [31:0] v482;
  wire signed [31:0] v483;
  wire signed [31:0] v484;
  wire signed [31:0] v485;
  wire signed [31:0] v486;
  wire signed [31:0] v487;
  wire signed [31:0] v488;
  wire signed [31:0] v489;
  wire signed [31:0] v490;
  wire signed [31:0] v491;
  wire signed [31:0] v492;
  wire signed [31:0] v493;
  wire signed [31:0] v494;
  wire signed [31:0] v495;
  wire signed [31:0] v496;
  wire signed [31:0] v497;
  wire signed [31:0] v498;
  wire signed [31:0] v499;
  wire signed [31:0] v500;
  wire signed [31:0] v501;
  wire signed [31:0] v502;
  wire signed [31:0] v503;
  wire signed [31:0] v504;
  wire signed [31:0] v505;
  wire signed [31:0] v506;
  wire signed [31:0] v507;
  wire signed [31:0] v508;
  wire signed [31:0] v509;
  wire signed [31:0] v510;
  wire signed [31:0] v511;
  wire signed [31:0] v512;
  wire signed [31:0] v513;
  wire signed [31:0] v514;
  wire signed [31:0] v515;
  wire signed [31:0] v516;
  wire signed [31:0] v517;
  wire signed [31:0] v518;
  wire signed [31:0] v519;
  wire signed [31:0] v520;
  wire signed [31:0] v521;
  wire signed [31:0] v522;
  wire signed [31:0] v523;
  wire signed [31:0] v524;
  wire signed [31:0] v525;
  wire signed [31:0] v526;
  wire signed [31:0] v527;
  wire signed [31:0] v528;
  wire signed [31:0] v529;
  wire signed [31:0] v530;
  wire signed [31:0] v531;
  wire signed [31:0] v532;
  wire signed [31:0] v533;
  wire signed [31:0] v534;
  wire signed [31:0] v535;
  wire signed [31:0] v536;
  wire signed [31:0] v537;
  wire signed [31:0] v538;
  wire signed [31:0] v539;
  wire signed [31:0] v540;
  wire signed [31:0] v541;
  wire signed [31:0] v542;
  wire signed [31:0] v543;
  wire signed [31:0] v544;
  wire signed [31:0] v545;
  wire signed [31:0] v546;
  wire signed [31:0] v547;
  wire signed [31:0] v548;
  wire signed [31:0] v549;
  wire signed [31:0] v550;
  wire signed [31:0] v551;
  wire signed [31:0] v552;
  wire signed [31:0] v553;
  wire signed [31:0] v554;
  wire signed [31:0] v555;
  wire signed [31:0] v556;
  wire signed [31:0] v557;
  wire signed [31:0] v558;
  wire signed [31:0] v559;
  wire signed [31:0] v560;
  wire signed [31:0] v561;
  wire signed [31:0] v562;
  wire signed [31:0] v563;
  wire signed [31:0] v564;
  wire signed [31:0] v565;
  wire signed [31:0] v566;
  wire signed [31:0] v567;
  wire signed [31:0] v568;
  wire signed [31:0] v569;
  wire signed [31:0] v570;
  wire signed [31:0] v571;
  wire signed [31:0] v572;
  wire signed [31:0] v573;
  wire signed [31:0] v574;
  wire signed [31:0] v575;
  wire signed [31:0] v576;
  wire signed [31:0] v577;
  wire signed [31:0] v578;
  wire signed [31:0] v579;
  wire signed [31:0] v580;
  wire signed [31:0] v581;
  wire signed [31:0] v582;
  wire signed [31:0] v583;
  wire signed [31:0] v584;
  wire signed [31:0] v585;
  wire signed [31:0] v586;
  wire signed [31:0] v587;
  wire signed [31:0] v588;
  wire signed [31:0] v589;
  wire signed [31:0] v590;
  wire signed [31:0] v591;
  wire signed [31:0] v592;
  wire signed [31:0] v593;
  wire signed [31:0] v594;
  wire signed [31:0] v595;
  wire signed [31:0] v596;
  wire signed [31:0] v597;
  wire signed [31:0] v598;
  wire signed [31:0] v599;
  wire signed [31:0] v600;
  wire signed [31:0] v601;
  wire signed [31:0] v602;
  wire signed [31:0] v603;
  wire signed [31:0] v604;
  wire signed [31:0] v605;
  wire signed [31:0] v606;
  wire signed [31:0] v607;
  wire signed [31:0] v608;
  wire signed [31:0] v609;
  wire signed [31:0] v610;
  wire signed [31:0] v611;
  wire signed [31:0] v612;
  wire signed [31:0] v613;
  wire signed [31:0] v614;
  wire signed [31:0] v615;
  wire signed [31:0] v616;
  wire signed [31:0] v617;
  wire signed [31:0] v618;
  wire signed [31:0] v619;
  wire signed [31:0] v620;
  wire signed [31:0] v621;
  wire signed [31:0] v622;
  wire signed [31:0] v623;
  wire signed [31:0] v624;
  wire signed [31:0] v625;
  wire signed [31:0] v626;
  wire signed [31:0] v627;
  wire signed [31:0] v628;
  wire signed [31:0] v629;
  wire signed [31:0] v630;
  wire signed [31:0] v631;
  wire signed [31:0] v632;
  wire signed [31:0] v633;
  wire signed [31:0] v634;
  wire signed [31:0] v635;
  wire signed [31:0] v636;
  wire signed [31:0] v637;
  wire signed [31:0] v638;
  wire signed [31:0] v639;
  wire signed [31:0] v640;
  wire signed [31:0] v641;
  wire signed [31:0] v642;
  wire signed [31:0] v643;
  wire signed [31:0] v644;
  wire signed [31:0] v645;
  wire signed [31:0] v646;
  wire signed [31:0] v647;
  wire signed [31:0] v648;
  wire signed [31:0] v649;
  wire signed [31:0] v650;
  wire signed [31:0] v651;
  wire signed [31:0] v652;
  wire signed [31:0] v653;
  wire signed [31:0] v654;
  wire signed [31:0] v655;
  wire signed [31:0] v656;
  wire signed [31:0] v657;
  wire signed [31:0] v658;
  wire signed [31:0] v659;
  wire signed [31:0] v660;
  wire signed [31:0] v661;
  wire signed [31:0] v662;
  wire signed [31:0] v663;
  wire signed [31:0] v664;
  wire signed [31:0] v665;
  wire signed [31:0] v666;
  wire signed [31:0] v667;
  wire signed [31:0] v668;
  wire signed [31:0] v669;
  wire signed [31:0] v670;
  wire signed [31:0] v671;
  wire signed [31:0] v672;
  wire signed [31:0] v673;
  wire signed [31:0] v674;
  wire signed [31:0] v675;
  wire signed [31:0] v676;
  wire signed [31:0] v677;
  wire signed [31:0] v678;
  wire signed [31:0] v679;
  wire signed [31:0] v680;
  wire signed [31:0] v681;
  wire signed [31:0] v682;
  wire signed [31:0] v683;
  wire signed [31:0] v684;
  wire signed [31:0] v685;
  wire signed [31:0] v686;
  wire signed [31:0] v687;
  wire signed [31:0] v688;
  wire signed [31:0] v689;
  wire signed [31:0] v690;
  wire signed [31:0] v691;
  wire signed [31:0] v692;
  wire signed [31:0] v693;
  wire signed [31:0] v694;
  wire signed [31:0] v695;
  wire signed [31:0] v696;
  wire signed [31:0] v697;
  wire signed [31:0] v698;
  wire signed [31:0] v699;
  wire signed [31:0] v700;
  wire signed [31:0] v701;
  wire signed [31:0] v702;
  wire signed [31:0] v703;
  wire signed [31:0] v704;
  wire signed [31:0] v705;
  wire signed [31:0] v706;
  wire signed [31:0] v707;
  wire signed [31:0] v708;
  wire signed [31:0] v709;
  wire signed [31:0] v710;
  wire signed [31:0] v711;
  wire signed [31:0] v712;
  wire signed [31:0] v713;
  wire signed [31:0] v714;
  wire signed [31:0] v715;
  wire signed [31:0] v716;
  wire signed [31:0] v717;
  wire signed [31:0] v718;
  wire signed [31:0] v719;
  wire signed [31:0] v720;
  wire signed [31:0] v721;
  wire signed [31:0] v722;
  wire signed [31:0] v723;
  wire signed [31:0] v724;
  wire signed [31:0] v725;
  wire signed [31:0] v726;
  wire signed [31:0] v727;
  wire signed [31:0] v728;
  wire signed [31:0] v729;
  wire signed [31:0] v730;
  wire signed [31:0] v731;
  wire signed [31:0] v732;
  wire signed [31:0] v733;
  wire signed [31:0] v734;
  wire signed [31:0] v735;
  wire signed [31:0] v736;
  wire signed [31:0] v737;
  wire signed [31:0] v738;
  wire signed [31:0] v739;
  wire signed [31:0] v740;
  wire signed [31:0] v741;
  wire signed [31:0] v742;
  wire signed [31:0] v743;
  wire signed [31:0] v744;
  wire signed [31:0] v745;
  wire signed [31:0] v746;
  wire signed [31:0] v747;
  wire signed [31:0] v748;
  wire signed [31:0] v749;
  wire signed [31:0] v750;
  wire signed [31:0] v751;
  wire signed [31:0] v752;
  wire signed [31:0] v753;
  wire signed [31:0] v754;
  wire signed [31:0] v755;
  wire signed [31:0] v756;
  wire signed [31:0] v757;
  wire signed [31:0] v758;
  wire signed [31:0] v759;
  wire signed [31:0] v760;
  wire signed [31:0] v761;
  wire signed [31:0] v762;
  wire signed [31:0] v763;
  wire signed [31:0] v764;
  wire signed [31:0] v765;
  wire signed [31:0] v766;
  wire signed [31:0] v767;
  wire signed [31:0] v768;
  wire signed [31:0] v769;
  wire signed [31:0] v770;
  wire signed [31:0] v771;
  wire signed [31:0] v772;
  wire signed [31:0] v773;
  wire signed [31:0] v774;
  wire signed [31:0] v775;
  wire signed [31:0] v776;
  wire signed [31:0] v777;
  wire signed [31:0] v778;
  wire signed [31:0] v779;
  wire signed [31:0] v780;
  wire signed [31:0] v781;
  wire signed [31:0] v782;
  wire signed [31:0] v783;
  wire signed [31:0] v784;
  wire signed [31:0] v785;
  wire signed [31:0] v786;
  wire signed [31:0] v787;
  wire signed [31:0] v788;
  wire signed [31:0] v789;
  wire signed [31:0] v790;
  wire signed [31:0] v791;
  wire signed [31:0] v792;
  wire signed [31:0] v793;
  wire signed [31:0] v794;
  wire signed [31:0] v795;
  wire signed [31:0] v796;
  wire signed [31:0] v797;
  wire signed [31:0] v798;
  wire signed [31:0] v799;
  wire signed [31:0] v800;
  wire signed [31:0] v801;
  wire signed [31:0] v802;
  wire signed [31:0] v803;
  wire signed [31:0] v804;
  wire signed [31:0] v805;
  wire signed [31:0] v806;
  wire signed [31:0] v807;
  wire signed [31:0] v808;
  wire signed [31:0] v809;
  wire signed [31:0] v810;
  wire signed [31:0] v811;
  wire signed [31:0] v812;
  wire signed [31:0] v813;
  wire signed [31:0] v814;
  wire signed [31:0] v815;
  wire signed [31:0] v816;
  wire signed [31:0] v817;
  wire signed [31:0] v818;
  wire signed [31:0] v819;
  wire signed [31:0] v820;
  wire signed [31:0] v821;
  wire signed [31:0] v822;
  wire signed [31:0] v823;
  wire signed [31:0] v824;
  wire signed [31:0] v825;
  wire signed [31:0] v826;
  wire signed [31:0] v827;
  wire signed [31:0] v828;
  wire signed [31:0] v829;
  wire signed [31:0] v830;
  wire signed [31:0] v831;
  wire signed [31:0] v832;
  wire signed [31:0] v833;
  wire signed [31:0] v834;
  wire signed [31:0] v835;
  wire signed [31:0] v836;
  wire signed [31:0] v837;
  wire signed [31:0] v838;
  wire signed [31:0] v839;
  wire signed [31:0] v840;
  wire signed [31:0] v841;
  wire signed [31:0] v842;
  wire signed [31:0] v843;
  wire signed [31:0] v844;
  wire signed [31:0] v845;
  wire signed [31:0] v846;
  wire signed [31:0] v847;
  wire signed [31:0] v848;
  wire signed [31:0] v849;
  wire signed [31:0] v850;
  wire signed [31:0] v851;
  wire signed [31:0] v852;
  wire signed [31:0] v853;
  wire signed [31:0] v854;
  wire signed [31:0] v855;
  wire signed [31:0] v856;
  wire signed [31:0] v857;
  wire signed [31:0] v858;
  wire signed [31:0] v859;
  wire signed [31:0] v860;
  wire signed [31:0] v861;
  wire signed [31:0] v862;
  wire signed [31:0] v863;
  wire signed [31:0] v864;
  wire signed [31:0] v865;
  wire signed [31:0] v866;
  wire signed [31:0] v867;
  wire signed [31:0] v868;
  wire signed [31:0] v869;
  wire signed [31:0] v870;
  wire signed [31:0] v871;
  wire signed [31:0] v872;
  wire signed [31:0] v873;
  wire signed [31:0] v874;
  wire signed [31:0] v875;
  wire signed [31:0] v876;
  wire signed [31:0] v877;
  wire signed [31:0] v878;
  wire signed [31:0] v879;
  wire signed [31:0] v880;
  wire signed [31:0] v881;
  wire signed [31:0] v882;
  wire signed [31:0] v883;
  wire signed [31:0] v884;
  wire signed [31:0] v885;
  wire signed [31:0] v886;
  wire signed [31:0] v887;
  wire signed [31:0] v888;
  wire signed [31:0] v889;
  wire signed [31:0] v890;
  wire signed [31:0] v891;
  wire signed [31:0] v892;
  wire signed [31:0] v893;
  wire signed [31:0] v894;
  wire signed [31:0] v895;
  wire signed [31:0] v896;
  wire signed [31:0] v897;
  wire signed [31:0] v898;
  wire signed [31:0] v899;
  wire signed [31:0] v900;
  wire signed [31:0] v901;
  wire signed [31:0] v902;
  wire signed [31:0] v903;
  wire signed [31:0] v904;
  wire signed [31:0] v905;
  wire signed [31:0] v906;
  wire signed [31:0] v907;
  wire signed [31:0] v908;
  wire signed [31:0] v909;
  wire signed [31:0] v910;
  wire signed [31:0] v911;
  wire signed [31:0] v912;
  wire signed [31:0] v913;
  wire signed [31:0] v914;
  wire signed [31:0] v915;
  wire signed [31:0] v916;
  wire signed [31:0] v917;
  wire signed [31:0] v918;
  wire signed [31:0] v919;
  wire signed [31:0] v920;
  wire signed [31:0] v921;
  wire signed [31:0] v922;
  wire signed [31:0] v923;
  wire signed [31:0] v924;
  wire signed [31:0] v925;
  wire signed [31:0] v926;
  wire signed [31:0] v927;
  wire signed [31:0] v928;
  wire signed [31:0] v929;
  wire signed [31:0] v930;
  wire signed [31:0] v931;
  wire signed [31:0] v932;
  wire signed [31:0] v933;
  wire signed [31:0] v934;
  wire signed [31:0] v935;
  wire signed [31:0] v936;
  wire signed [31:0] v937;
  wire signed [31:0] v938;
  wire signed [31:0] v939;
  wire signed [31:0] v940;
  wire signed [31:0] v941;
  wire signed [31:0] v942;
  wire signed [31:0] v943;
  wire signed [31:0] v944;
  wire signed [31:0] v945;
  wire signed [31:0] v946;
  wire signed [31:0] v947;
  wire signed [31:0] v948;
  wire signed [31:0] v949;
  wire signed [31:0] v950;
  wire signed [31:0] v951;
  wire signed [31:0] v952;
  wire signed [31:0] v953;
  wire signed [31:0] v954;
  wire signed [31:0] v955;
  wire signed [31:0] v956;
  wire signed [31:0] v957;
  wire signed [31:0] v958;
  wire signed [31:0] v959;
  wire signed [31:0] v960;
  wire signed [31:0] v961;
  wire signed [31:0] v962;
  wire signed [31:0] v963;
  wire signed [31:0] v964;
  wire signed [31:0] v965;
  wire signed [31:0] v966;
  wire signed [31:0] v967;
  wire signed [31:0] v968;
  wire signed [31:0] v969;
  wire signed [31:0] v970;
  wire signed [31:0] v971;
  wire signed [31:0] v972;
  wire signed [31:0] v973;
  wire signed [31:0] v974;
  wire signed [31:0] v975;
  wire signed [31:0] v976;
  wire signed [31:0] v977;
  wire signed [31:0] v978;
  wire signed [63:0] v979;
  wire signed [63:0] v980;
  wire signed [63:0] v981;
  wire v982;
  wire signed [63:0] v983;
  wire signed [63:0] v984;
  wire signed [63:0] v985;
  wire signed [31:0] v986;
  wire signed [31:0] v987;
  wire v988;
  wire signed [31:0] v989;
  wire v990;
  wire signed [31:0] v991;
  wire signed [7:0] v992;
  wire signed [63:0] v993;
  wire signed [63:0] v994;
  wire signed [63:0] v995;
  wire v996;
  wire signed [63:0] v997;
  wire signed [63:0] v998;
  wire signed [63:0] v999;
  wire signed [31:0] v1000;
  wire signed [31:0] v1001;
  wire v1002;
  wire signed [31:0] v1003;
  wire v1004;
  wire signed [31:0] v1005;
  wire signed [7:0] v1006;
  wire signed [63:0] v1007;
  wire signed [63:0] v1008;
  wire signed [63:0] v1009;
  wire v1010;
  wire signed [63:0] v1011;
  wire signed [63:0] v1012;
  wire signed [63:0] v1013;
  wire signed [31:0] v1014;
  wire signed [31:0] v1015;
  wire v1016;
  wire signed [31:0] v1017;
  wire v1018;
  wire signed [31:0] v1019;
  wire signed [7:0] v1020;
  wire signed [63:0] v1021;
  wire signed [63:0] v1022;
  wire signed [63:0] v1023;
  wire v1024;
  wire signed [63:0] v1025;
  wire signed [63:0] v1026;
  wire signed [63:0] v1027;
  wire signed [31:0] v1028;
  wire signed [31:0] v1029;
  wire v1030;
  wire signed [31:0] v1031;
  wire v1032;
  wire signed [31:0] v1033;
  wire signed [7:0] v1034;
  wire signed [63:0] v1035;
  wire signed [63:0] v1036;
  wire signed [63:0] v1037;
  wire v1038;
  wire signed [63:0] v1039;
  wire signed [63:0] v1040;
  wire signed [63:0] v1041;
  wire signed [31:0] v1042;
  wire signed [31:0] v1043;
  wire v1044;
  wire signed [31:0] v1045;
  wire v1046;
  wire signed [31:0] v1047;
  wire signed [7:0] v1048;
  wire signed [63:0] v1049;
  wire signed [63:0] v1050;
  wire signed [63:0] v1051;
  wire v1052;
  wire signed [63:0] v1053;
  wire signed [63:0] v1054;
  wire signed [63:0] v1055;
  wire signed [31:0] v1056;
  wire signed [31:0] v1057;
  wire v1058;
  wire signed [31:0] v1059;
  wire v1060;
  wire signed [31:0] v1061;
  wire signed [7:0] v1062;
  wire signed [63:0] v1063;
  wire signed [63:0] v1064;
  wire signed [63:0] v1065;
  wire v1066;
  wire signed [63:0] v1067;
  wire signed [63:0] v1068;
  wire signed [63:0] v1069;
  wire signed [31:0] v1070;
  wire signed [31:0] v1071;
  wire v1072;
  wire signed [31:0] v1073;
  wire v1074;
  wire signed [31:0] v1075;
  wire signed [7:0] v1076;
  wire signed [63:0] v1077;
  wire signed [63:0] v1078;
  wire signed [63:0] v1079;
  wire v1080;
  wire signed [63:0] v1081;
  wire signed [63:0] v1082;
  wire signed [63:0] v1083;
  wire signed [31:0] v1084;
  wire signed [31:0] v1085;
  wire v1086;
  wire signed [31:0] v1087;
  wire v1088;
  wire signed [31:0] v1089;
  wire signed [7:0] v1090;
  wire signed [63:0] v1091;
  wire signed [63:0] v1092;
  wire signed [63:0] v1093;
  wire v1094;
  wire signed [63:0] v1095;
  wire signed [63:0] v1096;
  wire signed [63:0] v1097;
  wire signed [31:0] v1098;
  wire signed [31:0] v1099;
  wire v1100;
  wire signed [31:0] v1101;
  wire v1102;
  wire signed [31:0] v1103;
  wire signed [7:0] v1104;
  wire signed [63:0] v1105;
  wire signed [63:0] v1106;
  wire signed [63:0] v1107;
  wire v1108;
  wire signed [63:0] v1109;
  wire signed [63:0] v1110;
  wire signed [63:0] v1111;
  wire signed [31:0] v1112;
  wire signed [31:0] v1113;
  wire v1114;
  wire signed [31:0] v1115;
  wire v1116;
  wire signed [31:0] v1117;
  wire signed [7:0] v1118;
  wire signed [63:0] v1119;
  wire signed [63:0] v1120;
  wire signed [63:0] v1121;
  wire v1122;
  wire signed [63:0] v1123;
  wire signed [63:0] v1124;
  wire signed [63:0] v1125;
  wire signed [31:0] v1126;
  wire signed [31:0] v1127;
  wire v1128;
  wire signed [31:0] v1129;
  wire v1130;
  wire signed [31:0] v1131;
  wire signed [7:0] v1132;
  wire signed [63:0] v1133;
  wire signed [63:0] v1134;
  wire signed [63:0] v1135;
  wire v1136;
  wire signed [63:0] v1137;
  wire signed [63:0] v1138;
  wire signed [63:0] v1139;
  wire signed [31:0] v1140;
  wire signed [31:0] v1141;
  wire v1142;
  wire signed [31:0] v1143;
  wire v1144;
  wire signed [31:0] v1145;
  wire signed [7:0] v1146;
  wire signed [63:0] v1147;
  wire signed [63:0] v1148;
  wire signed [63:0] v1149;
  wire v1150;
  wire signed [63:0] v1151;
  wire signed [63:0] v1152;
  wire signed [63:0] v1153;
  wire signed [31:0] v1154;
  wire signed [31:0] v1155;
  wire v1156;
  wire signed [31:0] v1157;
  wire v1158;
  wire signed [31:0] v1159;
  wire signed [7:0] v1160;
  wire signed [63:0] v1161;
  wire signed [63:0] v1162;
  wire signed [63:0] v1163;
  wire v1164;
  wire signed [63:0] v1165;
  wire signed [63:0] v1166;
  wire signed [63:0] v1167;
  wire signed [31:0] v1168;
  wire signed [31:0] v1169;
  wire v1170;
  wire signed [31:0] v1171;
  wire v1172;
  wire signed [31:0] v1173;
  wire signed [7:0] v1174;
  wire signed [63:0] v1175;
  wire signed [63:0] v1176;
  wire signed [63:0] v1177;
  wire v1178;
  wire signed [63:0] v1179;
  wire signed [63:0] v1180;
  wire signed [63:0] v1181;
  wire signed [31:0] v1182;
  wire signed [31:0] v1183;
  wire v1184;
  wire signed [31:0] v1185;
  wire v1186;
  wire signed [31:0] v1187;
  wire signed [7:0] v1188;
  wire signed [63:0] v1189;
  wire signed [63:0] v1190;
  wire signed [63:0] v1191;
  wire v1192;
  wire signed [63:0] v1193;
  wire signed [63:0] v1194;
  wire signed [63:0] v1195;
  wire signed [31:0] v1196;
  wire signed [31:0] v1197;
  wire v1198;
  wire signed [31:0] v1199;
  wire v1200;
  wire signed [31:0] v1201;
  wire signed [7:0] v1202;
  wire v1203;
  wire signed [7:0] v1204;
  wire v1205;
  wire signed [7:0] v1206;
  wire v1207;
  wire signed [7:0] v1208;
  wire v1209;
  wire signed [7:0] v1210;
  wire v1211;
  wire signed [7:0] v1212;
  wire v1213;
  wire signed [7:0] v1214;
  wire v1215;
  wire signed [7:0] v1216;
  wire v1217;
  wire signed [7:0] v1218;
  wire v1219;
  wire signed [7:0] v1220;
  wire v1221;
  wire signed [7:0] v1222;
  wire v1223;
  wire signed [7:0] v1224;
  wire v1225;
  wire signed [7:0] v1226;
  wire v1227;
  wire signed [7:0] v1228;
  wire v1229;
  wire signed [7:0] v1230;
  wire v1231;
  wire signed [7:0] v1232;
  wire v1233;
  wire signed [7:0] v1234;
  wire v1235;
  wire signed [7:0] v1236;
  wire v1237;
  wire signed [7:0] v1238;
  wire v1239;
  wire signed [7:0] v1240;
  wire v1241;
  wire signed [7:0] v1242;
  wire v1243;
  wire signed [7:0] v1244;
  wire v1245;
  wire signed [7:0] v1246;
  wire v1247;
  wire signed [7:0] v1248;
  wire v1249;
  wire signed [7:0] v1250;
  wire v1251;
  wire signed [7:0] v1252;
  wire v1253;
  wire signed [7:0] v1254;
  wire v1255;
  wire signed [7:0] v1256;
  wire v1257;
  wire signed [7:0] v1258;
  wire v1259;
  wire signed [7:0] v1260;
  wire v1261;
  wire signed [7:0] v1262;
  wire v1263;
  wire signed [7:0] v1264;
  wire v1265;
  wire signed [7:0] v1266;
  wire signed [31:0] v1267;
  wire signed [31:0] v1268;
  wire signed [31:0] v1269;
  wire signed [31:0] v1270;
  wire signed [31:0] v1271;
  wire signed [31:0] v1272;
  wire signed [31:0] v1273;
  wire signed [31:0] v1274;
  wire signed [31:0] v1275;
  wire signed [31:0] v1276;
  wire signed [31:0] v1277;
  wire signed [31:0] v1278;
  wire signed [31:0] v1279;
  wire signed [31:0] v1280;
  wire signed [31:0] v1281;
  wire signed [31:0] v1282;
  wire signed [31:0] v1283;
  wire signed [31:0] v1284;
  wire signed [31:0] v1285;
  wire signed [31:0] v1286;
  wire signed [31:0] v1287;
  wire signed [31:0] v1288;
  wire signed [31:0] v1289;
  wire signed [31:0] v1290;
  wire signed [31:0] v1291;
  wire signed [31:0] v1292;
  wire signed [31:0] v1293;
  wire signed [31:0] v1294;
  wire signed [31:0] v1295;
  wire signed [31:0] v1296;
  wire signed [31:0] v1297;
  wire signed [31:0] v1298;
  wire signed [31:0] v1299;
  wire signed [31:0] v1300;
  wire signed [31:0] v1301;
  wire signed [31:0] v1302;
  wire signed [31:0] v1303;
  wire signed [31:0] v1304;
  wire signed [31:0] v1305;
  wire signed [31:0] v1306;
  wire signed [31:0] v1307;
  wire signed [31:0] v1308;
  wire signed [31:0] v1309;
  wire signed [31:0] v1310;
  wire signed [31:0] v1311;
  wire signed [31:0] v1312;
  wire signed [31:0] v1313;
  wire signed [31:0] v1314;
  wire signed [31:0] v1315;
  wire signed [31:0] v1316;
  wire signed [31:0] v1317;
  wire signed [31:0] v1318;
  wire signed [31:0] v1319;
  wire signed [31:0] v1320;
  wire signed [31:0] v1321;
  wire signed [31:0] v1322;
  wire signed [31:0] v1323;
  wire signed [31:0] v1324;
  wire signed [31:0] v1325;
  wire signed [31:0] v1326;
  wire signed [31:0] v1327;
  wire signed [31:0] v1328;
  wire signed [31:0] v1329;
  wire signed [31:0] v1330;
  wire signed [63:0] v1331;
  wire signed [63:0] v1332;
  wire signed [63:0] v1333;
  wire v1334;
  wire signed [63:0] v1335;
  wire signed [63:0] v1336;
  wire signed [63:0] v1337;
  wire signed [31:0] v1338;
  wire signed [31:0] v1339;
  wire v1340;
  wire signed [31:0] v1341;
  wire v1342;
  wire signed [31:0] v1343;
  wire signed [7:0] v1344;

  assign v2 = 0;
  assign v3 = -128;
  assign v4 = 1073741824;
  assign v5 = -1073741824;
  assign v6 = 127;
  assign v7 = -128;
  assign v8 = 127;
  assign v9 = 5;
  assign v10 = 36;
  assign v11 = 1630361836;
  assign v12 = 34359738368;
  assign v13 = 37;
  assign v14 = 1561796795;
  assign v15 = 68719476736;
  assign v16 = 38;
  assign v17 = 137438953472;
  assign v18 = 2039655736;
  assign v19 = 429;
  assign v20 = -729;
  assign v21 = 1954;
  assign v22 = 610;
  assign v23 = 241;
  assign v24 = -471;
  assign v25 = -35;
  assign v26 = -867;
  assign v27 = 571;
  assign v28 = 581;
  assign v29 = 4260;
  assign v30 = 3943;
  assign v31 = 591;
  assign v32 = -889;
  assign v33 = -5103;
  assign v34 = -5438;
  assign v35 = -5515;
  assign v36 = -1352;
  assign v37 = -1500;
  assign v38 = -4152;
  assign v39 = -84;
  assign v40 = 3396;
  assign v41 = 1981;
  assign v42 = -5581;
  assign v43 = -6964;
  assign v44 = 3407;
  assign v45 = -7217;
  assign v46 = -9;
  assign v47 = -54;
  assign v48 = 57;
  assign v49 = 71;
  assign v50 = 104;
  assign v51 = 115;
  assign v52 = 98;
  assign v53 = 99;
  assign v54 = 64;
  assign v55 = -26;
  assign v56 = 25;
  assign v57 = -82;
  assign v58 = 68;
  assign v59 = 95;
  assign v60 = 86;
  assign v61 = -12;
  assign v62 = 26;
  assign v63 = -19;
  assign v64 = 9;
  assign v65 = 33;
  assign v66 = 36;
  assign v67 = -32;
  assign v68 = -17;
  assign v69 = -68;
  assign v70 = -11;
  assign v71 = -6;
  assign v72 = 3;
  assign v73 = -36;
  assign v74 = -46;
  assign v75 = 2;
  assign v76 = 6;
  assign v77 = -7;
  assign v78 = -15;
  assign v79 = -45;
  assign v80 = 39;
  assign v81 = -31;
  assign v82 = -5;
  assign v83 = -21;
  assign v84 = -37;
  assign v85 = -28;
  assign v86 = 23;
  assign v87 = -4;
  assign v88 = 18;
  assign v89 = 21;
  assign v90 = 30;
  assign v91 = 16;
  assign v92 = -2;
  assign v93 = 20;
  assign v94 = -38;
  assign v95 = 28;
  assign v96 = -8;
  assign v97 = -13;
  assign v98 = -30;
  assign v99 = -29;
  assign v100 = -23;
  assign v101 = 7;
  assign v102 = 11;
  assign v103 = 4;
  assign v104 = 27;
  assign v105 = -34;
  assign v106 = -20;
  assign v107 = 35;
  assign v108 = 10;
  assign v109 = 34;
  assign v110 = -64;
  assign v111 = 17;
  assign v112 = 12;
  assign v113 = -27;
  assign v114 = -24;
  assign v115 = -3;
  assign v116 = 38;
  assign v117 = -25;
  assign v118 = -22;
  assign v119 = 37;
  assign v120 = 29;
  assign v121 = 32;
  assign v122 = 55;
  assign v123 = 22;
  assign v124 = 24;
  assign v125 = 46;
  assign v126 = -39;
  assign v127 = -40;
  assign v128 = 19;
  assign v129 = -60;
  assign v130 = 13;
  assign v131 = -42;
  assign v132 = 31;
  assign v133 = -41;
  assign v134 = -58;
  assign v135 = 62;
  assign v136 = -57;
  assign v137 = 8;
  assign v138 = 15;
  assign v139 = -18;
  assign v140 = 41;
  assign v141 = 88;
  assign v142 = 59;
  assign v143 = -59;
  assign v144 = {{24{arg1[7]}}, arg1};
  assign v145 = v144 - v3;
  assign v146 = v145 * v46;
  assign v147 = v145 * v47;
  assign v148 = v145 * v48;
  assign v149 = v145 * v49;
  assign v150 = v145 * v50;
  assign v151 = v145 * v51;
  assign v152 = v145 * v52;
  assign v153 = v145 * v53;
  assign v154 = v145 * v54;
  assign v155 = v145 * v55;
  assign v156 = v145 * v6;
  assign v157 = v145 * v56;
  assign v158 = v145 * v57;
  assign v159 = v145 * v58;
  assign v160 = v145 * v59;
  assign v161 = v145 * v60;
  assign v162 = v148 + v34;
  assign v163 = v149 + v35;
  assign v164 = v150 + v36;
  assign v165 = v151 + v37;
  assign v166 = v152 + v38;
  assign v167 = v153 + v39;
  assign v168 = v154 + v40;
  assign v169 = v156 + v41;
  assign v170 = v157 + v42;
  assign v171 = v159 + v43;
  assign v172 = v160 + v44;
  assign v173 = v161 + v45;
  assign v174 = {{32{v146[31]}}, v146};
  assign v175 = v174 * v18;
  assign v176 = v175 + v17;
  assign v177 = v146 >= v2;
  assign v178 = v177 ? v4 : v5;
  assign v179 = v178 + v176;
  assign v180 = v179 >>> v16;
  assign v181 = v180[31:0];
  assign v182 = v181 + v3;
  assign v183 = v182 < v3;
  assign v184 = v183 ? v3 : v182;
  assign v185 = v182 > v6;
  assign v186 = v185 ? v6 : v184;
  assign v187 = v186[7:0];
  assign v188 = {{32{v147[31]}}, v147};
  assign v189 = v188 * v18;
  assign v190 = v189 + v17;
  assign v191 = v147 >= v2;
  assign v192 = v191 ? v4 : v5;
  assign v193 = v192 + v190;
  assign v194 = v193 >>> v16;
  assign v195 = v194[31:0];
  assign v196 = v195 + v3;
  assign v197 = v196 < v3;
  assign v198 = v197 ? v3 : v196;
  assign v199 = v196 > v6;
  assign v200 = v199 ? v6 : v198;
  assign v201 = v200[7:0];
  assign v202 = {{32{v162[31]}}, v162};
  assign v203 = v202 * v18;
  assign v204 = v203 + v17;
  assign v205 = v162 >= v2;
  assign v206 = v205 ? v4 : v5;
  assign v207 = v206 + v204;
  assign v208 = v207 >>> v16;
  assign v209 = v208[31:0];
  assign v210 = v209 + v3;
  assign v211 = v210 < v3;
  assign v212 = v211 ? v3 : v210;
  assign v213 = v210 > v6;
  assign v214 = v213 ? v6 : v212;
  assign v215 = v214[7:0];
  assign v216 = {{32{v163[31]}}, v163};
  assign v217 = v216 * v18;
  assign v218 = v217 + v17;
  assign v219 = v163 >= v2;
  assign v220 = v219 ? v4 : v5;
  assign v221 = v220 + v218;
  assign v222 = v221 >>> v16;
  assign v223 = v222[31:0];
  assign v224 = v223 + v3;
  assign v225 = v224 < v3;
  assign v226 = v225 ? v3 : v224;
  assign v227 = v224 > v6;
  assign v228 = v227 ? v6 : v226;
  assign v229 = v228[7:0];
  assign v230 = {{32{v164[31]}}, v164};
  assign v231 = v230 * v18;
  assign v232 = v231 + v17;
  assign v233 = v164 >= v2;
  assign v234 = v233 ? v4 : v5;
  assign v235 = v234 + v232;
  assign v236 = v235 >>> v16;
  assign v237 = v236[31:0];
  assign v238 = v237 + v3;
  assign v239 = v238 < v3;
  assign v240 = v239 ? v3 : v238;
  assign v241 = v238 > v6;
  assign v242 = v241 ? v6 : v240;
  assign v243 = v242[7:0];
  assign v244 = {{32{v165[31]}}, v165};
  assign v245 = v244 * v18;
  assign v246 = v245 + v17;
  assign v247 = v165 >= v2;
  assign v248 = v247 ? v4 : v5;
  assign v249 = v248 + v246;
  assign v250 = v249 >>> v16;
  assign v251 = v250[31:0];
  assign v252 = v251 + v3;
  assign v253 = v252 < v3;
  assign v254 = v253 ? v3 : v252;
  assign v255 = v252 > v6;
  assign v256 = v255 ? v6 : v254;
  assign v257 = v256[7:0];
  assign v258 = {{32{v166[31]}}, v166};
  assign v259 = v258 * v18;
  assign v260 = v259 + v17;
  assign v261 = v166 >= v2;
  assign v262 = v261 ? v4 : v5;
  assign v263 = v262 + v260;
  assign v264 = v263 >>> v16;
  assign v265 = v264[31:0];
  assign v266 = v265 + v3;
  assign v267 = v266 < v3;
  assign v268 = v267 ? v3 : v266;
  assign v269 = v266 > v6;
  assign v270 = v269 ? v6 : v268;
  assign v271 = v270[7:0];
  assign v272 = {{32{v167[31]}}, v167};
  assign v273 = v272 * v18;
  assign v274 = v273 + v17;
  assign v275 = v167 >= v2;
  assign v276 = v275 ? v4 : v5;
  assign v277 = v276 + v274;
  assign v278 = v277 >>> v16;
  assign v279 = v278[31:0];
  assign v280 = v279 + v3;
  assign v281 = v280 < v3;
  assign v282 = v281 ? v3 : v280;
  assign v283 = v280 > v6;
  assign v284 = v283 ? v6 : v282;
  assign v285 = v284[7:0];
  assign v286 = {{32{v168[31]}}, v168};
  assign v287 = v286 * v18;
  assign v288 = v287 + v17;
  assign v289 = v168 >= v2;
  assign v290 = v289 ? v4 : v5;
  assign v291 = v290 + v288;
  assign v292 = v291 >>> v16;
  assign v293 = v292[31:0];
  assign v294 = v293 + v3;
  assign v295 = v294 < v3;
  assign v296 = v295 ? v3 : v294;
  assign v297 = v294 > v6;
  assign v298 = v297 ? v6 : v296;
  assign v299 = v298[7:0];
  assign v300 = {{32{v155[31]}}, v155};
  assign v301 = v300 * v18;
  assign v302 = v301 + v17;
  assign v303 = v155 >= v2;
  assign v304 = v303 ? v4 : v5;
  assign v305 = v304 + v302;
  assign v306 = v305 >>> v16;
  assign v307 = v306[31:0];
  assign v308 = v307 + v3;
  assign v309 = v308 < v3;
  assign v310 = v309 ? v3 : v308;
  assign v311 = v308 > v6;
  assign v312 = v311 ? v6 : v310;
  assign v313 = v312[7:0];
  assign v314 = {{32{v169[31]}}, v169};
  assign v315 = v314 * v18;
  assign v316 = v315 + v17;
  assign v317 = v169 >= v2;
  assign v318 = v317 ? v4 : v5;
  assign v319 = v318 + v316;
  assign v320 = v319 >>> v16;
  assign v321 = v320[31:0];
  assign v322 = v321 + v3;
  assign v323 = v322 < v3;
  assign v324 = v323 ? v3 : v322;
  assign v325 = v322 > v6;
  assign v326 = v325 ? v6 : v324;
  assign v327 = v326[7:0];
  assign v328 = {{32{v170[31]}}, v170};
  assign v329 = v328 * v18;
  assign v330 = v329 + v17;
  assign v331 = v170 >= v2;
  assign v332 = v331 ? v4 : v5;
  assign v333 = v332 + v330;
  assign v334 = v333 >>> v16;
  assign v335 = v334[31:0];
  assign v336 = v335 + v3;
  assign v337 = v336 < v3;
  assign v338 = v337 ? v3 : v336;
  assign v339 = v336 > v6;
  assign v340 = v339 ? v6 : v338;
  assign v341 = v340[7:0];
  assign v342 = {{32{v158[31]}}, v158};
  assign v343 = v342 * v18;
  assign v344 = v343 + v17;
  assign v345 = v158 >= v2;
  assign v346 = v345 ? v4 : v5;
  assign v347 = v346 + v344;
  assign v348 = v347 >>> v16;
  assign v349 = v348[31:0];
  assign v350 = v349 + v3;
  assign v351 = v350 < v3;
  assign v352 = v351 ? v3 : v350;
  assign v353 = v350 > v6;
  assign v354 = v353 ? v6 : v352;
  assign v355 = v354[7:0];
  assign v356 = {{32{v171[31]}}, v171};
  assign v357 = v356 * v18;
  assign v358 = v357 + v17;
  assign v359 = v171 >= v2;
  assign v360 = v359 ? v4 : v5;
  assign v361 = v360 + v358;
  assign v362 = v361 >>> v16;
  assign v363 = v362[31:0];
  assign v364 = v363 + v3;
  assign v365 = v364 < v3;
  assign v366 = v365 ? v3 : v364;
  assign v367 = v364 > v6;
  assign v368 = v367 ? v6 : v366;
  assign v369 = v368[7:0];
  assign v370 = {{32{v172[31]}}, v172};
  assign v371 = v370 * v18;
  assign v372 = v371 + v17;
  assign v373 = v172 >= v2;
  assign v374 = v373 ? v4 : v5;
  assign v375 = v374 + v372;
  assign v376 = v375 >>> v16;
  assign v377 = v376[31:0];
  assign v378 = v377 + v3;
  assign v379 = v378 < v3;
  assign v380 = v379 ? v3 : v378;
  assign v381 = v378 > v6;
  assign v382 = v381 ? v6 : v380;
  assign v383 = v382[7:0];
  assign v384 = {{32{v173[31]}}, v173};
  assign v385 = v384 * v18;
  assign v386 = v385 + v17;
  assign v387 = v173 >= v2;
  assign v388 = v387 ? v4 : v5;
  assign v389 = v388 + v386;
  assign v390 = v389 >>> v16;
  assign v391 = v390[31:0];
  assign v392 = v391 + v3;
  assign v393 = v392 < v3;
  assign v394 = v393 ? v3 : v392;
  assign v395 = v392 > v6;
  assign v396 = v395 ? v6 : v394;
  assign v397 = v396[7:0];
  assign v398 = v187 < v7;
  assign v399 = v398 ? v7 : v187;
  assign v400 = v187 > v8;
  assign v401 = v400 ? v8 : v399;
  assign v402 = v201 < v7;
  assign v403 = v402 ? v7 : v201;
  assign v404 = v201 > v8;
  assign v405 = v404 ? v8 : v403;
  assign v406 = v215 < v7;
  assign v407 = v406 ? v7 : v215;
  assign v408 = v215 > v8;
  assign v409 = v408 ? v8 : v407;
  assign v410 = v229 < v7;
  assign v411 = v410 ? v7 : v229;
  assign v412 = v229 > v8;
  assign v413 = v412 ? v8 : v411;
  assign v414 = v243 < v7;
  assign v415 = v414 ? v7 : v243;
  assign v416 = v243 > v8;
  assign v417 = v416 ? v8 : v415;
  assign v418 = v257 < v7;
  assign v419 = v418 ? v7 : v257;
  assign v420 = v257 > v8;
  assign v421 = v420 ? v8 : v419;
  assign v422 = v271 < v7;
  assign v423 = v422 ? v7 : v271;
  assign v424 = v271 > v8;
  assign v425 = v424 ? v8 : v423;
  assign v426 = v285 < v7;
  assign v427 = v426 ? v7 : v285;
  assign v428 = v285 > v8;
  assign v429 = v428 ? v8 : v427;
  assign v430 = v299 < v7;
  assign v431 = v430 ? v7 : v299;
  assign v432 = v299 > v8;
  assign v433 = v432 ? v8 : v431;
  assign v434 = v313 < v7;
  assign v435 = v434 ? v7 : v313;
  assign v436 = v313 > v8;
  assign v437 = v436 ? v8 : v435;
  assign v438 = v327 < v7;
  assign v439 = v438 ? v7 : v327;
  assign v440 = v327 > v8;
  assign v441 = v440 ? v8 : v439;
  assign v442 = v341 < v7;
  assign v443 = v442 ? v7 : v341;
  assign v444 = v341 > v8;
  assign v445 = v444 ? v8 : v443;
  assign v446 = v355 < v7;
  assign v447 = v446 ? v7 : v355;
  assign v448 = v355 > v8;
  assign v449 = v448 ? v8 : v447;
  assign v450 = v369 < v7;
  assign v451 = v450 ? v7 : v369;
  assign v452 = v369 > v8;
  assign v453 = v452 ? v8 : v451;
  assign v454 = v383 < v7;
  assign v455 = v454 ? v7 : v383;
  assign v456 = v383 > v8;
  assign v457 = v456 ? v8 : v455;
  assign v458 = v397 < v7;
  assign v459 = v458 ? v7 : v397;
  assign v460 = v397 > v8;
  assign v461 = v460 ? v8 : v459;
  assign v462 = {{24{v401[7]}}, v401};
  assign v463 = v462 - v3;
  assign v464 = v463 * v61;
  assign v465 = {{24{v405[7]}}, v405};
  assign v466 = v465 - v3;
  assign v467 = v466 * v62;
  assign v468 = v464 + v467;
  assign v469 = {{24{v409[7]}}, v409};
  assign v470 = v469 - v3;
  assign v471 = v470 * v63;
  assign v472 = v468 + v471;
  assign v473 = {{24{v413[7]}}, v413};
  assign v474 = v473 - v3;
  assign v475 = v474 * v64;
  assign v476 = v472 + v475;
  assign v477 = {{24{v417[7]}}, v417};
  assign v478 = v477 - v3;
  assign v479 = v478 * v56;
  assign v480 = v476 + v479;
  assign v481 = {{24{v421[7]}}, v421};
  assign v482 = v481 - v3;
  assign v483 = v482 * v65;
  assign v484 = v480 + v483;
  assign v485 = {{24{v425[7]}}, v425};
  assign v486 = v485 - v3;
  assign v487 = v486 * v61;
  assign v488 = v484 + v487;
  assign v489 = {{24{v429[7]}}, v429};
  assign v490 = v489 - v3;
  assign v491 = v490 * v66;
  assign v492 = v488 + v491;
  assign v493 = {{24{v433[7]}}, v433};
  assign v494 = v493 - v3;
  assign v495 = v494 * v67;
  assign v496 = v492 + v495;
  assign v497 = {{24{v437[7]}}, v437};
  assign v498 = v497 - v3;
  assign v499 = v498 * v65;
  assign v500 = v496 + v499;
  assign v501 = {{24{v441[7]}}, v441};
  assign v502 = v501 - v3;
  assign v503 = v502 * v68;
  assign v504 = v500 + v503;
  assign v505 = {{24{v445[7]}}, v445};
  assign v506 = v505 - v3;
  assign v507 = v506 * v69;
  assign v508 = v504 + v507;
  assign v509 = {{24{v449[7]}}, v449};
  assign v510 = v509 - v3;
  assign v511 = v510 * v46;
  assign v512 = v508 + v511;
  assign v513 = {{24{v453[7]}}, v453};
  assign v514 = v513 - v3;
  assign v515 = v514 * v70;
  assign v516 = v512 + v515;
  assign v517 = {{24{v457[7]}}, v457};
  assign v518 = v517 - v3;
  assign v519 = v518 * v71;
  assign v520 = v516 + v519;
  assign v521 = {{24{v461[7]}}, v461};
  assign v522 = v521 - v3;
  assign v523 = v522 * v56;
  assign v524 = v520 + v523;
  assign v525 = v463 * v72;
  assign v526 = v466 * v73;
  assign v527 = v525 + v526;
  assign v528 = v470 * v74;
  assign v529 = v527 + v528;
  assign v530 = v474 * v75;
  assign v531 = v529 + v530;
  assign v532 = v478 * v76;
  assign v533 = v531 + v532;
  assign v534 = v482 * v77;
  assign v535 = v533 + v534;
  assign v536 = v535 + v487;
  assign v537 = v490 * v75;
  assign v538 = v536 + v537;
  assign v539 = v538 - v494;
  assign v540 = v498 * v71;
  assign v541 = v539 + v540;
  assign v542 = v541 + v503;
  assign v543 = v506 * v78;
  assign v544 = v542 + v543;
  assign v545 = v510 * v68;
  assign v546 = v544 + v545;
  assign v547 = v514 * v79;
  assign v548 = v546 + v547;
  assign v549 = v518 * v80;
  assign v550 = v548 + v549;
  assign v551 = v522 * v81;
  assign v552 = v550 + v551;
  assign v553 = v463 * v82;
  assign v554 = v466 * v80;
  assign v555 = v553 + v554;
  assign v556 = v470 * v25;
  assign v557 = v555 + v556;
  assign v558 = v474 * v83;
  assign v559 = v557 + v558;
  assign v560 = v478 * v84;
  assign v561 = v559 + v560;
  assign v562 = v482 * v85;
  assign v563 = v561 + v562;
  assign v564 = v486 * v9;
  assign v565 = v563 + v564;
  assign v566 = v490 * v62;
  assign v567 = v565 + v566;
  assign v568 = v494 * v86;
  assign v569 = v567 + v568;
  assign v570 = v498 * v87;
  assign v571 = v569 + v570;
  assign v572 = v502 * v66;
  assign v573 = v571 + v572;
  assign v574 = v506 * v88;
  assign v575 = v573 + v574;
  assign v576 = v510 * v89;
  assign v577 = v575 + v576;
  assign v578 = v514 * v68;
  assign v579 = v577 + v578;
  assign v580 = v518 * v90;
  assign v581 = v579 + v580;
  assign v582 = v522 * v85;
  assign v583 = v581 + v582;
  assign v584 = v463 * v91;
  assign v585 = v466 * v92;
  assign v586 = v584 + v585;
  assign v587 = v470 * v93;
  assign v588 = v586 + v587;
  assign v589 = v474 * v94;
  assign v590 = v588 + v589;
  assign v591 = v478 * v95;
  assign v592 = v590 + v591;
  assign v593 = v482 * v96;
  assign v594 = v592 + v593;
  assign v595 = v486 * v97;
  assign v596 = v594 + v595;
  assign v597 = v490 * v78;
  assign v598 = v596 + v597;
  assign v599 = v494 * v68;
  assign v600 = v598 + v599;
  assign v601 = v498 * v98;
  assign v602 = v600 + v601;
  assign v603 = v502 * v97;
  assign v604 = v602 + v603;
  assign v605 = v506 * v64;
  assign v606 = v604 + v605;
  assign v607 = v510 * v99;
  assign v608 = v606 + v607;
  assign v609 = v514 * v100;
  assign v610 = v608 + v609;
  assign v611 = v518 * v63;
  assign v612 = v610 + v611;
  assign v613 = v522 * v99;
  assign v614 = v612 + v613;
  assign v615 = v463 * v85;
  assign v616 = v466 * v89;
  assign v617 = v615 + v616;
  assign v618 = v470 * v101;
  assign v619 = v617 + v618;
  assign v620 = v474 * v102;
  assign v621 = v619 + v620;
  assign v622 = v478 * v103;
  assign v623 = v621 + v622;
  assign v624 = v482 * v104;
  assign v625 = v623 + v624;
  assign v626 = v486 * v62;
  assign v627 = v625 + v626;
  assign v628 = v490 * v92;
  assign v629 = v627 + v628;
  assign v630 = v494 * v83;
  assign v631 = v629 + v630;
  assign v632 = v631 + v498;
  assign v633 = v502 * v105;
  assign v634 = v632 + v633;
  assign v635 = v506 * v65;
  assign v636 = v634 + v635;
  assign v637 = v510 * v55;
  assign v638 = v636 + v637;
  assign v639 = v514 * v102;
  assign v640 = v638 + v639;
  assign v641 = v518 * v106;
  assign v642 = v640 + v641;
  assign v643 = v522 * v72;
  assign v644 = v642 + v643;
  assign v645 = v463 * v107;
  assign v646 = v466 * v108;
  assign v647 = v645 + v646;
  assign v648 = v470 * v109;
  assign v649 = v647 + v648;
  assign v650 = v474 * v66;
  assign v651 = v649 + v650;
  assign v652 = v478 * v90;
  assign v653 = v651 + v652;
  assign v654 = v482 * v80;
  assign v655 = v653 + v654;
  assign v656 = v486 * v72;
  assign v657 = v655 + v656;
  assign v658 = v490 * v55;
  assign v659 = v657 + v658;
  assign v660 = v494 * v72;
  assign v661 = v659 + v660;
  assign v662 = v498 * v66;
  assign v663 = v661 + v662;
  assign v664 = v663 - v502;
  assign v665 = v506 * v110;
  assign v666 = v664 + v665;
  assign v667 = v510 * v111;
  assign v668 = v666 + v667;
  assign v669 = v514 * v96;
  assign v670 = v668 + v669;
  assign v671 = v518 * v87;
  assign v672 = v670 + v671;
  assign v673 = v522 * v78;
  assign v674 = v672 + v673;
  assign v675 = v463 * v111;
  assign v676 = v466 * v112;
  assign v677 = v675 + v676;
  assign v678 = v470 * v70;
  assign v679 = v677 + v678;
  assign v680 = v474 * v67;
  assign v681 = v679 + v680;
  assign v682 = v478 * v97;
  assign v683 = v681 + v682;
  assign v684 = v482 * v101;
  assign v685 = v683 + v684;
  assign v686 = v486 * v86;
  assign v687 = v685 + v686;
  assign v688 = v490 * v113;
  assign v689 = v687 + v688;
  assign v690 = v494 * v114;
  assign v691 = v689 + v690;
  assign v692 = v498 * v63;
  assign v693 = v691 + v692;
  assign v694 = v502 * v71;
  assign v695 = v693 + v694;
  assign v696 = v506 * v73;
  assign v697 = v695 + v696;
  assign v698 = v510 * v114;
  assign v699 = v697 + v698;
  assign v700 = v514 * v107;
  assign v701 = v699 + v700;
  assign v702 = v518 * v82;
  assign v703 = v701 + v702;
  assign v704 = v522 * v101;
  assign v705 = v703 + v704;
  assign v706 = v463 * v25;
  assign v707 = v466 * v82;
  assign v708 = v706 + v707;
  assign v709 = v470 * v115;
  assign v710 = v708 + v709;
  assign v711 = v478 * v93;
  assign v712 = v710 + v711;
  assign v713 = v482 * v116;
  assign v714 = v712 + v713;
  assign v715 = v486 * v111;
  assign v716 = v714 + v715;
  assign v717 = v490 * v86;
  assign v718 = v716 + v717;
  assign v719 = v494 * v117;
  assign v720 = v718 + v719;
  assign v721 = v498 * v78;
  assign v722 = v720 + v721;
  assign v723 = v502 * v111;
  assign v724 = v722 + v723;
  assign v725 = v506 * v118;
  assign v726 = v724 + v725;
  assign v727 = v510 * v75;
  assign v728 = v726 + v727;
  assign v729 = v514 * v116;
  assign v730 = v728 + v729;
  assign v731 = v518 * v103;
  assign v732 = v730 + v731;
  assign v733 = v522 * v103;
  assign v734 = v732 + v733;
  assign v735 = v463 * v119;
  assign v736 = v466 * v65;
  assign v737 = v735 + v736;
  assign v738 = v470 * v120;
  assign v739 = v737 + v738;
  assign v740 = v474 * v108;
  assign v741 = v739 + v740;
  assign v742 = v741 + v560;
  assign v743 = v482 * v120;
  assign v744 = v742 + v743;
  assign v745 = v486 * v73;
  assign v746 = v744 + v745;
  assign v747 = v490 * v121;
  assign v748 = v746 + v747;
  assign v749 = v748 + v494;
  assign v750 = v749 + v540;
  assign v751 = v502 * v99;
  assign v752 = v750 + v751;
  assign v753 = v506 * v122;
  assign v754 = v752 + v753;
  assign v755 = v510 * v102;
  assign v756 = v754 + v755;
  assign v757 = v514 * v78;
  assign v758 = v756 + v757;
  assign v759 = v518 * v62;
  assign v760 = v758 + v759;
  assign v761 = v522 * v123;
  assign v762 = v760 + v761;
  assign v763 = v463 * v68;
  assign v764 = v466 * v95;
  assign v765 = v763 + v764;
  assign v766 = v470 * v117;
  assign v767 = v765 + v766;
  assign v768 = v474 * v72;
  assign v769 = v767 + v768;
  assign v770 = v478 * v67;
  assign v771 = v769 + v770;
  assign v772 = v482 * v123;
  assign v773 = v771 + v772;
  assign v774 = v486 * v75;
  assign v775 = v773 + v774;
  assign v776 = v490 * v72;
  assign v777 = v775 + v776;
  assign v778 = v494 * v65;
  assign v779 = v777 + v778;
  assign v780 = v498 * v124;
  assign v781 = v779 + v780;
  assign v782 = v502 * v64;
  assign v783 = v781 + v782;
  assign v784 = v506 * v125;
  assign v785 = v783 + v784;
  assign v786 = v510 * v126;
  assign v787 = v785 + v786;
  assign v788 = v514 * v113;
  assign v789 = v787 + v788;
  assign v790 = v518 * v93;
  assign v791 = v789 + v790;
  assign v792 = v522 * v102;
  assign v793 = v791 + v792;
  assign v794 = v463 * v118;
  assign v795 = v794 + v467;
  assign v796 = v470 * v87;
  assign v797 = v795 + v796;
  assign v798 = v474 * v127;
  assign v799 = v797 + v798;
  assign v800 = v478 * v128;
  assign v801 = v799 + v800;
  assign v802 = v486 * v129;
  assign v803 = v801 + v802;
  assign v804 = v490 * v127;
  assign v805 = v803 + v804;
  assign v806 = v494 * v106;
  assign v807 = v805 + v806;
  assign v808 = v498 * v126;
  assign v809 = v807 + v808;
  assign v810 = v502 * v92;
  assign v811 = v809 + v810;
  assign v812 = v506 * v130;
  assign v813 = v811 + v812;
  assign v814 = v510 * v56;
  assign v815 = v813 + v814;
  assign v816 = v514 * v121;
  assign v817 = v815 + v816;
  assign v818 = v518 * v127;
  assign v819 = v817 + v818;
  assign v820 = v522 * v131;
  assign v821 = v819 + v820;
  assign v822 = v463 * v98;
  assign v823 = v466 * v132;
  assign v824 = v822 + v823;
  assign v825 = v470 * v100;
  assign v826 = v824 + v825;
  assign v827 = v474 * v133;
  assign v828 = v826 + v827;
  assign v829 = v478 * v47;
  assign v830 = v828 + v829;
  assign v831 = v482 * v98;
  assign v832 = v830 + v831;
  assign v833 = v486 * v25;
  assign v834 = v832 + v833;
  assign v835 = v490 * v134;
  assign v836 = v834 + v835;
  assign v837 = v494 * v128;
  assign v838 = v836 + v837;
  assign v839 = v498 * v117;
  assign v840 = v838 + v839;
  assign v841 = v502 * v103;
  assign v842 = v840 + v841;
  assign v843 = v506 * v135;
  assign v844 = v842 + v843;
  assign v845 = v844 + v514;
  assign v846 = v845 + v790;
  assign v847 = v522 * v136;
  assign v848 = v846 + v847;
  assign v849 = v463 * v84;
  assign v850 = v466 * v117;
  assign v851 = v849 + v850;
  assign v852 = v470 * v89;
  assign v853 = v851 + v852;
  assign v854 = v474 * v89;
  assign v855 = v853 + v854;
  assign v856 = v478 * v70;
  assign v857 = v855 + v856;
  assign v858 = v482 * v76;
  assign v859 = v857 + v858;
  assign v860 = v486 * v131;
  assign v861 = v859 + v860;
  assign v862 = v861 + v566;
  assign v863 = v494 * v73;
  assign v864 = v862 + v863;
  assign v865 = v498 * v64;
  assign v866 = v864 + v865;
  assign v867 = v502 * v109;
  assign v868 = v866 + v867;
  assign v869 = v506 * v92;
  assign v870 = v868 + v869;
  assign v871 = v510 * v137;
  assign v872 = v870 + v871;
  assign v873 = v514 * v75;
  assign v874 = v872 + v873;
  assign v875 = v518 * v128;
  assign v876 = v874 + v875;
  assign v877 = v522 * v68;
  assign v878 = v876 + v877;
  assign v879 = v463 * v56;
  assign v880 = v466 * v90;
  assign v881 = v879 + v880;
  assign v882 = v470 * v98;
  assign v883 = v881 + v882;
  assign v884 = v883 + v475;
  assign v885 = v478 * v115;
  assign v886 = v884 + v885;
  assign v887 = v482 * v97;
  assign v888 = v886 + v887;
  assign v889 = v486 * v93;
  assign v890 = v888 + v889;
  assign v891 = v490 * v25;
  assign v892 = v890 + v891;
  assign v893 = v494 * v94;
  assign v894 = v892 + v893;
  assign v895 = v498 * v121;
  assign v896 = v894 + v895;
  assign v897 = v502 * v126;
  assign v898 = v896 + v897;
  assign v899 = v506 * v138;
  assign v900 = v898 + v899;
  assign v901 = v900 + v607;
  assign v902 = v514 * v77;
  assign v903 = v901 + v902;
  assign v904 = v518 * v46;
  assign v905 = v903 + v904;
  assign v906 = v522 * v139;
  assign v907 = v905 + v906;
  assign v908 = v463 * v100;
  assign v909 = v466 * v66;
  assign v910 = v908 + v909;
  assign v911 = v470 * v55;
  assign v912 = v910 + v911;
  assign v913 = v474 * v140;
  assign v914 = v912 + v913;
  assign v915 = v914 + v684;
  assign v916 = v486 * v123;
  assign v917 = v915 + v916;
  assign v918 = v490 * v98;
  assign v919 = v917 + v918;
  assign v920 = v494 * v90;
  assign v921 = v919 + v920;
  assign v922 = v498 * v130;
  assign v923 = v921 + v922;
  assign v924 = v502 * v107;
  assign v925 = v923 + v924;
  assign v926 = v506 * v79;
  assign v927 = v925 + v926;
  assign v928 = v510 * v25;
  assign v929 = v927 + v928;
  assign v930 = v514 * v46;
  assign v931 = v929 + v930;
  assign v932 = v931 + v790;
  assign v933 = v522 * v71;
  assign v934 = v932 + v933;
  assign v935 = v463 * v137;
  assign v936 = v466 * v109;
  assign v937 = v935 + v936;
  assign v938 = v470 * v116;
  assign v939 = v937 + v938;
  assign v940 = v474 * v65;
  assign v941 = v939 + v940;
  assign v942 = v478 * v64;
  assign v943 = v941 + v942;
  assign v944 = v482 * v137;
  assign v945 = v943 + v944;
  assign v946 = v486 * v138;
  assign v947 = v945 + v946;
  assign v948 = v490 * v102;
  assign v949 = v947 + v948;
  assign v950 = v949 + v495;
  assign v951 = v498 * v88;
  assign v952 = v950 + v951;
  assign v953 = v502 * v61;
  assign v954 = v952 + v953;
  assign v955 = v506 * v6;
  assign v956 = v954 + v955;
  assign v957 = v510 * v73;
  assign v958 = v956 + v957;
  assign v959 = v514 * v141;
  assign v960 = v958 + v959;
  assign v961 = v518 * v113;
  assign v962 = v960 + v961;
  assign v963 = v522 * v116;
  assign v964 = v962 + v963;
  assign v965 = v524 + v20;
  assign v966 = v552 + v21;
  assign v967 = v583 + v22;
  assign v968 = v644 + v23;
  assign v969 = v674 + v24;
  assign v970 = v705 + v25;
  assign v971 = v734 + v26;
  assign v972 = v762 + v27;
  assign v973 = v793 + v28;
  assign v974 = v821 + v29;
  assign v975 = v848 + v30;
  assign v976 = v878 + v31;
  assign v977 = v934 + v32;
  assign v978 = v964 + v33;
  assign v979 = {{32{v965[31]}}, v965};
  assign v980 = v979 * v14;
  assign v981 = v980 + v15;
  assign v982 = v965 >= v2;
  assign v983 = v982 ? v4 : v5;
  assign v984 = v983 + v981;
  assign v985 = v984 >>> v13;
  assign v986 = v985[31:0];
  assign v987 = v986 + v3;
  assign v988 = v987 < v3;
  assign v989 = v988 ? v3 : v987;
  assign v990 = v987 > v6;
  assign v991 = v990 ? v6 : v989;
  assign v992 = v991[7:0];
  assign v993 = {{32{v966[31]}}, v966};
  assign v994 = v993 * v14;
  assign v995 = v994 + v15;
  assign v996 = v966 >= v2;
  assign v997 = v996 ? v4 : v5;
  assign v998 = v997 + v995;
  assign v999 = v998 >>> v13;
  assign v1000 = v999[31:0];
  assign v1001 = v1000 + v3;
  assign v1002 = v1001 < v3;
  assign v1003 = v1002 ? v3 : v1001;
  assign v1004 = v1001 > v6;
  assign v1005 = v1004 ? v6 : v1003;
  assign v1006 = v1005[7:0];
  assign v1007 = {{32{v967[31]}}, v967};
  assign v1008 = v1007 * v14;
  assign v1009 = v1008 + v15;
  assign v1010 = v967 >= v2;
  assign v1011 = v1010 ? v4 : v5;
  assign v1012 = v1011 + v1009;
  assign v1013 = v1012 >>> v13;
  assign v1014 = v1013[31:0];
  assign v1015 = v1014 + v3;
  assign v1016 = v1015 < v3;
  assign v1017 = v1016 ? v3 : v1015;
  assign v1018 = v1015 > v6;
  assign v1019 = v1018 ? v6 : v1017;
  assign v1020 = v1019[7:0];
  assign v1021 = {{32{v614[31]}}, v614};
  assign v1022 = v1021 * v14;
  assign v1023 = v1022 + v15;
  assign v1024 = v614 >= v2;
  assign v1025 = v1024 ? v4 : v5;
  assign v1026 = v1025 + v1023;
  assign v1027 = v1026 >>> v13;
  assign v1028 = v1027[31:0];
  assign v1029 = v1028 + v3;
  assign v1030 = v1029 < v3;
  assign v1031 = v1030 ? v3 : v1029;
  assign v1032 = v1029 > v6;
  assign v1033 = v1032 ? v6 : v1031;
  assign v1034 = v1033[7:0];
  assign v1035 = {{32{v968[31]}}, v968};
  assign v1036 = v1035 * v14;
  assign v1037 = v1036 + v15;
  assign v1038 = v968 >= v2;
  assign v1039 = v1038 ? v4 : v5;
  assign v1040 = v1039 + v1037;
  assign v1041 = v1040 >>> v13;
  assign v1042 = v1041[31:0];
  assign v1043 = v1042 + v3;
  assign v1044 = v1043 < v3;
  assign v1045 = v1044 ? v3 : v1043;
  assign v1046 = v1043 > v6;
  assign v1047 = v1046 ? v6 : v1045;
  assign v1048 = v1047[7:0];
  assign v1049 = {{32{v969[31]}}, v969};
  assign v1050 = v1049 * v14;
  assign v1051 = v1050 + v15;
  assign v1052 = v969 >= v2;
  assign v1053 = v1052 ? v4 : v5;
  assign v1054 = v1053 + v1051;
  assign v1055 = v1054 >>> v13;
  assign v1056 = v1055[31:0];
  assign v1057 = v1056 + v3;
  assign v1058 = v1057 < v3;
  assign v1059 = v1058 ? v3 : v1057;
  assign v1060 = v1057 > v6;
  assign v1061 = v1060 ? v6 : v1059;
  assign v1062 = v1061[7:0];
  assign v1063 = {{32{v970[31]}}, v970};
  assign v1064 = v1063 * v14;
  assign v1065 = v1064 + v15;
  assign v1066 = v970 >= v2;
  assign v1067 = v1066 ? v4 : v5;
  assign v1068 = v1067 + v1065;
  assign v1069 = v1068 >>> v13;
  assign v1070 = v1069[31:0];
  assign v1071 = v1070 + v3;
  assign v1072 = v1071 < v3;
  assign v1073 = v1072 ? v3 : v1071;
  assign v1074 = v1071 > v6;
  assign v1075 = v1074 ? v6 : v1073;
  assign v1076 = v1075[7:0];
  assign v1077 = {{32{v971[31]}}, v971};
  assign v1078 = v1077 * v14;
  assign v1079 = v1078 + v15;
  assign v1080 = v971 >= v2;
  assign v1081 = v1080 ? v4 : v5;
  assign v1082 = v1081 + v1079;
  assign v1083 = v1082 >>> v13;
  assign v1084 = v1083[31:0];
  assign v1085 = v1084 + v3;
  assign v1086 = v1085 < v3;
  assign v1087 = v1086 ? v3 : v1085;
  assign v1088 = v1085 > v6;
  assign v1089 = v1088 ? v6 : v1087;
  assign v1090 = v1089[7:0];
  assign v1091 = {{32{v972[31]}}, v972};
  assign v1092 = v1091 * v14;
  assign v1093 = v1092 + v15;
  assign v1094 = v972 >= v2;
  assign v1095 = v1094 ? v4 : v5;
  assign v1096 = v1095 + v1093;
  assign v1097 = v1096 >>> v13;
  assign v1098 = v1097[31:0];
  assign v1099 = v1098 + v3;
  assign v1100 = v1099 < v3;
  assign v1101 = v1100 ? v3 : v1099;
  assign v1102 = v1099 > v6;
  assign v1103 = v1102 ? v6 : v1101;
  assign v1104 = v1103[7:0];
  assign v1105 = {{32{v973[31]}}, v973};
  assign v1106 = v1105 * v14;
  assign v1107 = v1106 + v15;
  assign v1108 = v973 >= v2;
  assign v1109 = v1108 ? v4 : v5;
  assign v1110 = v1109 + v1107;
  assign v1111 = v1110 >>> v13;
  assign v1112 = v1111[31:0];
  assign v1113 = v1112 + v3;
  assign v1114 = v1113 < v3;
  assign v1115 = v1114 ? v3 : v1113;
  assign v1116 = v1113 > v6;
  assign v1117 = v1116 ? v6 : v1115;
  assign v1118 = v1117[7:0];
  assign v1119 = {{32{v974[31]}}, v974};
  assign v1120 = v1119 * v14;
  assign v1121 = v1120 + v15;
  assign v1122 = v974 >= v2;
  assign v1123 = v1122 ? v4 : v5;
  assign v1124 = v1123 + v1121;
  assign v1125 = v1124 >>> v13;
  assign v1126 = v1125[31:0];
  assign v1127 = v1126 + v3;
  assign v1128 = v1127 < v3;
  assign v1129 = v1128 ? v3 : v1127;
  assign v1130 = v1127 > v6;
  assign v1131 = v1130 ? v6 : v1129;
  assign v1132 = v1131[7:0];
  assign v1133 = {{32{v975[31]}}, v975};
  assign v1134 = v1133 * v14;
  assign v1135 = v1134 + v15;
  assign v1136 = v975 >= v2;
  assign v1137 = v1136 ? v4 : v5;
  assign v1138 = v1137 + v1135;
  assign v1139 = v1138 >>> v13;
  assign v1140 = v1139[31:0];
  assign v1141 = v1140 + v3;
  assign v1142 = v1141 < v3;
  assign v1143 = v1142 ? v3 : v1141;
  assign v1144 = v1141 > v6;
  assign v1145 = v1144 ? v6 : v1143;
  assign v1146 = v1145[7:0];
  assign v1147 = {{32{v976[31]}}, v976};
  assign v1148 = v1147 * v14;
  assign v1149 = v1148 + v15;
  assign v1150 = v976 >= v2;
  assign v1151 = v1150 ? v4 : v5;
  assign v1152 = v1151 + v1149;
  assign v1153 = v1152 >>> v13;
  assign v1154 = v1153[31:0];
  assign v1155 = v1154 + v3;
  assign v1156 = v1155 < v3;
  assign v1157 = v1156 ? v3 : v1155;
  assign v1158 = v1155 > v6;
  assign v1159 = v1158 ? v6 : v1157;
  assign v1160 = v1159[7:0];
  assign v1161 = {{32{v907[31]}}, v907};
  assign v1162 = v1161 * v14;
  assign v1163 = v1162 + v15;
  assign v1164 = v907 >= v2;
  assign v1165 = v1164 ? v4 : v5;
  assign v1166 = v1165 + v1163;
  assign v1167 = v1166 >>> v13;
  assign v1168 = v1167[31:0];
  assign v1169 = v1168 + v3;
  assign v1170 = v1169 < v3;
  assign v1171 = v1170 ? v3 : v1169;
  assign v1172 = v1169 > v6;
  assign v1173 = v1172 ? v6 : v1171;
  assign v1174 = v1173[7:0];
  assign v1175 = {{32{v977[31]}}, v977};
  assign v1176 = v1175 * v14;
  assign v1177 = v1176 + v15;
  assign v1178 = v977 >= v2;
  assign v1179 = v1178 ? v4 : v5;
  assign v1180 = v1179 + v1177;
  assign v1181 = v1180 >>> v13;
  assign v1182 = v1181[31:0];
  assign v1183 = v1182 + v3;
  assign v1184 = v1183 < v3;
  assign v1185 = v1184 ? v3 : v1183;
  assign v1186 = v1183 > v6;
  assign v1187 = v1186 ? v6 : v1185;
  assign v1188 = v1187[7:0];
  assign v1189 = {{32{v978[31]}}, v978};
  assign v1190 = v1189 * v14;
  assign v1191 = v1190 + v15;
  assign v1192 = v978 >= v2;
  assign v1193 = v1192 ? v4 : v5;
  assign v1194 = v1193 + v1191;
  assign v1195 = v1194 >>> v13;
  assign v1196 = v1195[31:0];
  assign v1197 = v1196 + v3;
  assign v1198 = v1197 < v3;
  assign v1199 = v1198 ? v3 : v1197;
  assign v1200 = v1197 > v6;
  assign v1201 = v1200 ? v6 : v1199;
  assign v1202 = v1201[7:0];
  assign v1203 = v992 < v7;
  assign v1204 = v1203 ? v7 : v992;
  assign v1205 = v992 > v8;
  assign v1206 = v1205 ? v8 : v1204;
  assign v1207 = v1006 < v7;
  assign v1208 = v1207 ? v7 : v1006;
  assign v1209 = v1006 > v8;
  assign v1210 = v1209 ? v8 : v1208;
  assign v1211 = v1020 < v7;
  assign v1212 = v1211 ? v7 : v1020;
  assign v1213 = v1020 > v8;
  assign v1214 = v1213 ? v8 : v1212;
  assign v1215 = v1034 < v7;
  assign v1216 = v1215 ? v7 : v1034;
  assign v1217 = v1034 > v8;
  assign v1218 = v1217 ? v8 : v1216;
  assign v1219 = v1048 < v7;
  assign v1220 = v1219 ? v7 : v1048;
  assign v1221 = v1048 > v8;
  assign v1222 = v1221 ? v8 : v1220;
  assign v1223 = v1062 < v7;
  assign v1224 = v1223 ? v7 : v1062;
  assign v1225 = v1062 > v8;
  assign v1226 = v1225 ? v8 : v1224;
  assign v1227 = v1076 < v7;
  assign v1228 = v1227 ? v7 : v1076;
  assign v1229 = v1076 > v8;
  assign v1230 = v1229 ? v8 : v1228;
  assign v1231 = v1090 < v7;
  assign v1232 = v1231 ? v7 : v1090;
  assign v1233 = v1090 > v8;
  assign v1234 = v1233 ? v8 : v1232;
  assign v1235 = v1104 < v7;
  assign v1236 = v1235 ? v7 : v1104;
  assign v1237 = v1104 > v8;
  assign v1238 = v1237 ? v8 : v1236;
  assign v1239 = v1118 < v7;
  assign v1240 = v1239 ? v7 : v1118;
  assign v1241 = v1118 > v8;
  assign v1242 = v1241 ? v8 : v1240;
  assign v1243 = v1132 < v7;
  assign v1244 = v1243 ? v7 : v1132;
  assign v1245 = v1132 > v8;
  assign v1246 = v1245 ? v8 : v1244;
  assign v1247 = v1146 < v7;
  assign v1248 = v1247 ? v7 : v1146;
  assign v1249 = v1146 > v8;
  assign v1250 = v1249 ? v8 : v1248;
  assign v1251 = v1160 < v7;
  assign v1252 = v1251 ? v7 : v1160;
  assign v1253 = v1160 > v8;
  assign v1254 = v1253 ? v8 : v1252;
  assign v1255 = v1174 < v7;
  assign v1256 = v1255 ? v7 : v1174;
  assign v1257 = v1174 > v8;
  assign v1258 = v1257 ? v8 : v1256;
  assign v1259 = v1188 < v7;
  assign v1260 = v1259 ? v7 : v1188;
  assign v1261 = v1188 > v8;
  assign v1262 = v1261 ? v8 : v1260;
  assign v1263 = v1202 < v7;
  assign v1264 = v1263 ? v7 : v1202;
  assign v1265 = v1202 > v8;
  assign v1266 = v1265 ? v8 : v1264;
  assign v1267 = {{24{v1206[7]}}, v1206};
  assign v1268 = v1267 - v3;
  assign v1269 = v1268 * v126;
  assign v1270 = {{24{v1210[7]}}, v1210};
  assign v1271 = v1270 - v3;
  assign v1272 = v1271 * v142;
  assign v1273 = v1269 + v1272;
  assign v1274 = {{24{v1214[7]}}, v1214};
  assign v1275 = v1274 - v3;
  assign v1276 = v1275 * v80;
  assign v1277 = v1273 + v1276;
  assign v1278 = {{24{v1218[7]}}, v1218};
  assign v1279 = v1278 - v3;
  assign v1280 = v1279 * v89;
  assign v1281 = v1277 + v1280;
  assign v1282 = {{24{v1222[7]}}, v1222};
  assign v1283 = v1282 - v3;
  assign v1284 = v1283 * v95;
  assign v1285 = v1281 + v1284;
  assign v1286 = {{24{v1226[7]}}, v1226};
  assign v1287 = v1286 - v3;
  assign v1288 = v1287 * v67;
  assign v1289 = v1285 + v1288;
  assign v1290 = {{24{v1230[7]}}, v1230};
  assign v1291 = v1290 - v3;
  assign v1292 = v1291 * v105;
  assign v1293 = v1289 + v1292;
  assign v1294 = {{24{v1234[7]}}, v1234};
  assign v1295 = v1294 - v3;
  assign v1296 = v1295 * v25;
  assign v1297 = v1293 + v1296;
  assign v1298 = {{24{v1238[7]}}, v1238};
  assign v1299 = v1298 - v3;
  assign v1300 = v1299 * v138;
  assign v1301 = v1297 + v1300;
  assign v1302 = {{24{v1242[7]}}, v1242};
  assign v1303 = v1302 - v3;
  assign v1304 = v1303 * v104;
  assign v1305 = v1301 + v1304;
  assign v1306 = {{24{v1246[7]}}, v1246};
  assign v1307 = v1306 - v3;
  assign v1308 = v1307 * v143;
  assign v1309 = v1305 + v1308;
  assign v1310 = {{24{v1250[7]}}, v1250};
  assign v1311 = v1310 - v3;
  assign v1312 = v1311 * v133;
  assign v1313 = v1309 + v1312;
  assign v1314 = {{24{v1254[7]}}, v1254};
  assign v1315 = v1314 - v3;
  assign v1316 = v1315 * v88;
  assign v1317 = v1313 + v1316;
  assign v1318 = {{24{v1258[7]}}, v1258};
  assign v1319 = v1318 - v3;
  assign v1320 = v1319 * v25;
  assign v1321 = v1317 + v1320;
  assign v1322 = {{24{v1262[7]}}, v1262};
  assign v1323 = v1322 - v3;
  assign v1324 = v1323 * v77;
  assign v1325 = v1321 + v1324;
  assign v1326 = {{24{v1266[7]}}, v1266};
  assign v1327 = v1326 - v3;
  assign v1328 = v1327 * v6;
  assign v1329 = v1325 + v1328;
  assign v1330 = v1329 + v19;
  assign v1331 = {{32{v1330[31]}}, v1330};
  assign v1332 = v1331 * v11;
  assign v1333 = v1332 + v12;
  assign v1334 = v1330 >= v2;
  assign v1335 = v1334 ? v4 : v5;
  assign v1336 = v1335 + v1333;
  assign v1337 = v1336 >>> v10;
  assign v1338 = v1337[31:0];
  assign v1339 = v1338 + v9;
  assign v1340 = v1339 < v3;
  assign v1341 = v1340 ? v3 : v1339;
  assign v1342 = v1339 > v6;
  assign v1343 = v1342 ? v6 : v1341;
  assign v1344 = v1343[7:0];
  assign _out_ = v1344;
endmodule
